* NMOS Id-Vd

.include nmos.modelcard
.option abstol=1e-12
.option gmin=0

* Define parameterization for tests
.param
+ v_gate=1.2
+ v_drain=1.2
+ v_bulk=0.0
+ NF=1

* Define voltage sources, set to appropriate parameter values
vg gate  0 'v_gate'
vd drain 0 'v_drain'
vs bulk  0 'v_bulk'

m1 drain gate 0 bulk n1 W=10.0u L=0.09u NF='NF'
